`timescale 1ns / 1ps


module s12(
    input logic [31:0] a,
    output logic [31:0] y
    );
    // sal by 2
    assign y = {a[29:0], 2'b00};

endmodule
